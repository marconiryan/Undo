module main

pub fn asd() {
	println('asd')
}
