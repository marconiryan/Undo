module log

pub fn parse(){
	println('pasrse')
}
